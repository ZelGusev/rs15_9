public static void MakePowTable(uint New_GF_Byte_poly, uint New_GF_Byte_prim_memb, bool ShowMessageboxes) {
	//Если есть функция умножения, то составить таблицу степеней и логарифмов
	//не составляет никакого труда, ведь возведение в степень – есть умножение
	//несколько раз подряд
	//Здесь создаётся таблица степеней методом последовательного умножения
	//примитивного члена (как правило выбирают число 2, но здесь это может
	//быть любое число).
	//Затем таблица проверяется на наличие повторяющихся значений. Если нет
	//повторяющихся значений, то выбранный примитивный член и порождающий
	//полином сохраняются вместе с вычисленными таблицами.
	//для параметра New_GF_Byte_prim_memb валидны следующие значения:
	//285, 299, 301, 333, 351, 355, 357, 361, 369, 391, 397, 425, 251, 463,
	//487, 501.
	
	//Этот массив можно сделать на единицу меньше, так как для поля GF[256]
	//верно, что a^0= ^255, но чтобы не путаться оставляю 256 элементов массива.
	byte[] tmp_GF_256_power_a = new byte[256];	
	byte[] tmp_GF_256_log_a = new byte[256];
	GF_256_power_a = new byte[256];
	GF_256_log_a = new byte[256];

	uint tmp_GF_Byte_poly = New_GF_Byte_poly;
	uint tmp_GF_Byte_prim_memb = New_GF_Byte_prim_memb;

	//Пропишем тривиальные вещи как то: a^0=1 и a^1=a, и наоборот
	tmp_GF_256_power_a[0] = 1; 
	tmp_GF_256_log_a[1] = 0;
	tmp_GF_256_power_a[1] = (byte)tmp_GF_Byte_prim_memb;
	tmp_GF_256_log_a[tmp_GF_Byte_prim_memb] = 1;
	//Остальные члены поля
	for (int i = 2; i < 256; i++) {
		tmp_GF_256_power_a[i] = (byte)GF_b2_Aryth.Galois_b2_ext_mult(tmp_GF_Byte_prim_memb, tmp_GF_256_power_a[i - 1], tmp_GF_Byte_poly);
	//Для значения степени "0" тут проходят 2 значения: 1 и 255. Это надо учесть
		if(0 != tmp_GF_256_power_a[i]) {
			tmp_GF_256_log_a[tmp_GF_256_power_a[i]] = (byte)i;
		}
	}

	bool Ok = true;
	//Для поля GF[256] верно, что a^0 = a^255. Так что проверка
	//не затрагивает степень 255
	for (int i = 0; i <= 254; i++) {
		for (int j = 0; j <= 254; j++) {
			if (i != j) {
				if (tmp_GF_256_power_a[i] == tmp_GF_256_power_a[j]) {
					Ok = false;
				}
			}
		}
	}

	//Копируем в используемые таблицы, если нет повторов в таблице
	//степеней выбранного примитивного члена
	if (Ok) {
		for (int i = 0; i < 256; i++) {
			GF_256_power_a[i] = tmp_GF_256_power_a[i];
		}
		for (int i = 0; i < 256; i++) {
			GF_256_log_a[i] = tmp_GF_256_log_a[i];
		}
		GF_256_poly = tmp_GF_Byte_poly;
		GF_256_prim_memb = tmp_GF_Byte_prim_memb;
		if (ShowMessageboxes) { MessageBox.Show("Всё хорошо. При таком сочетании порождающего полинома и примитивного члена в таблице степеней примитивного члена (a^1 .. a^255) нет повторений."); }
	} else {
		if (ShowMessageboxes) { MessageBox.Show("Всё плохо! При таком сочетании порождающего полинома и примитивного члена в таблице степеней примитивного члена есть повторяющиеся значения."); }
	}
}

public static byte Pow_a(int Degr) {
	//Возведение примитивного члена в степень. Свойство степени в поле 
	//Галуа GF[256] таково, что степень примитивного члена 0 равна
	//степени 255; 1 - 256; 2 - 527 и так далее.
	if (0 <= Degr && Degr < 255) {
		return GF_256_power_a[Degr];
	} else {
		int TmpDegr = Glob.IntMod(Degr);
		TmpDegr %= 255; 
		//Хоть и не существует отрицательных чисел в поле Галуа, здесь под
		//отрицательной степенью подразумевается число обратное.
		if (Degr < 0) {
			TmpDegr = 255 - TmpDegr;
		}
		return GF_256_power_a[TmpDegr];
	}
}

public static byte Log_a(byte Arg) {
	//Логарифм по основанию примитивного члена
	if (0 == Arg) {
		throw new Exception("Argument cannot be zero in GF_Byte.Log_a(Arg)");		
	//Логарифм единицы в GF[256] равен нулю и 255, так как a^0==a^255.
	//Для кодирования Рида-Соломона выбираем 0.
	} else if (1 == Arg) { 
		return 0;
	}else {
		return GF_256_log_a[Arg];
	}
}

public static byte Inverse(byte Arg) {
	//Можно обойтись и без этой функции и писать Div(1, Arg)
	if (1 == Arg) { return 1; }
	return GF_256_power_a[255 - GF_256_log_a[Arg]];
}

public static byte Add(byte a1, byte a2) {
	//Сложение таково же как и вычитание - побитовое "ИЛИ"
	return (byte)(a1 ^ a2);
}

public static byte Sub(byte s1, byte s2) {
	//Вычитание таково же как и сложение - побитовое "ИЛИ"
	return (byte)(s1 ^ s2);
}

public static byte Mult(byte m1, byte m2) {
	//Умножение с использованием таблиц степеней и логарифмов.
	//Довольно таки быстрая операция
	if (0 == m1 || 0 == m2) { return 0; }
	return Pow_a(Log_a(m1) + Log_a(m2));
}

public static byte Div(byte d1, byte d2) {
	//Деление с использованием таблиц степеней и логарифмов.
	if (0 == d2) { throw new Exception("Division by zero"); }
	if (0 == d1) { return 0; }
	return Pow_a(Log_a(d1) - Log_a(d2));
}

public static byte Pow(byte b, int p) {
	//Возведение в степень с помощью таблиц логарифмов и степеней.
	 //Так как нуль в степени нуль равно одному, сначала проверяем
	 //на равенство нулю показателя
	if (0 == p) { return 1; }
	if (0 == b) { return 0; }
	byte BaseLog = GF_256_log_a[b];            
	int TmpDegr = Glob.IntMod(p);
	TmpDegr = TmpDegr * BaseLog;
	TmpDegr %= 255;
	if (p < 0) {
		TmpDegr = 255 - TmpDegr;
	}
	return GF_256_power_a[(byte)TmpDegr];}

module gf2_8_mul(
        input wire [7:0]    A   ,  //被乘数
        input wire [7:0]    B   ,  //乘数
        
        output wire[7:0]    P      //积
    );
    
    //多项式幂次为7的两个数相乘展开后最高幂次为14,对应15bit二进制数
    //超出GF(2^8)表示范围,先暂存,后续进行处理
    wire [14:0]  t_reg       ;   
    
    //依据伽罗华域GF(2^8)中的运算规则,预处理多项式的每一位
    assign t_reg[0]  = (A[0] & B[0]); 
    assign t_reg[1]  = (A[0] & B[1]) ^ (A[1] & B[0]);
    assign t_reg[2]  = (A[0] & B[2]) ^ (A[1] & B[1]) ^ (A[2] & B[0]);
    assign t_reg[3]  = (A[0] & B[3]) ^ (A[1] & B[2]) ^ (A[2] & B[1]) ^ (A[3] & B[0]);
    assign t_reg[4]  = (A[0] & B[4]) ^ (A[1] & B[3]) ^ (A[2] & B[2]) ^ (A[3] & B[1]) ^ (A[4] & B[0]);
    assign t_reg[5]  = (A[0] & B[5]) ^ (A[1] & B[4]) ^ (A[2] & B[3]) ^ (A[3] & B[2]) ^ (A[4] & B[1]) ^ (A[5] & B[0]); 
    assign t_reg[6]  = (A[0] & B[6]) ^ (A[1] & B[5]) ^ (A[2] & B[4]) ^ (A[3] & B[3]) ^ (A[4] & B[2]) ^ (A[5] & B[1]) ^ (A[6] & B[0]);
    assign t_reg[7]  = (A[0] & B[7]) ^ (A[1] & B[6]) ^ (A[2] & B[5]) ^ (A[3] & B[4]) ^ (A[4] & B[3]) ^ (A[5] & B[2]) ^ (A[6] & B[1]) ^ (A[7] & B[0]);
    assign t_reg[8]  = (A[1] & B[7]) ^ (A[2] & B[6]) ^ (A[3] & B[5]) ^ (A[4] & B[4]) ^ (A[5] & B[3]) ^ (A[6] & B[2]) ^ (A[7] & B[1]);
    assign t_reg[9]  = (A[2] & B[7]) ^ (A[3] & B[6]) ^ (A[4] & B[5]) ^ (A[5] & B[4]) ^ (A[6] & B[3]) ^ (A[7] & B[2]);
    assign t_reg[10] = (A[3] & B[7]) ^ (A[4] & B[6]) ^ (A[5] & B[5]) ^ (A[6] & B[4]) ^ (A[7] & B[3]);
    assign t_reg[11] = (A[4] & B[7]) ^ (A[5] & B[6]) ^ (A[6] & B[5]) ^ (A[7] & B[4]);
    assign t_reg[12] = (A[5] & B[7]) ^ (A[6] & B[6]) ^ (A[7] & B[5]);
    assign t_reg[13] = (A[6] & B[7]) ^ (A[7] & B[6]);
    assign t_reg[14] = (A[7] & B[7]);
    
    
    assign P[0] = t_reg[0] ^ t_reg[8]  ^ t_reg[12] ^ t_reg[13] ^ t_reg[14];
    assign P[1] = t_reg[1] ^ t_reg[9]  ^ t_reg[13] ^ t_reg[14]            ;
    assign P[2] = t_reg[2] ^ t_reg[8]  ^ t_reg[10] ^ t_reg[12] ^ t_reg[13];
    assign P[3] = t_reg[3] ^ t_reg[8]  ^ t_reg[9]  ^ t_reg[11] ^ t_reg[12];
    assign P[4] = t_reg[4] ^ t_reg[8]  ^ t_reg[9]  ^ t_reg[10] ^ t_reg[14];
    assign P[5] = t_reg[5] ^ t_reg[9]  ^ t_reg[10] ^ t_reg[11]            ;
    assign P[6] = t_reg[6] ^ t_reg[10] ^ t_reg[11] ^ t_reg[12]            ;
    assign P[7] = t_reg[7] ^ t_reg[11] ^ t_reg[12] ^ t_reg[13]            ;
    
endmodule

    GF(2^2) x^2+x+1
GF(2^3) x^3+x+1
GF(2^4) x^4+x+1
GF(2^5) x^5+x^2+1
GF(2^6) x^6+x+1
GF(2^7) x^7+x^3+1
GF(2^8) x^8+x^4+x^3+x^2+1
GF(2^9) x^9+x^4+1
GF(2^10) x^10+x^3+1
GF(2^11) x^11+x^2+1
GF(2^12) x^12+x^6+x^4+x+1
GF(2^13) x^13+x^4+x^3+x+1
GF(2^14) x^14+x^10+x^6+x+1
GF(2^15) x^15+x+1
GF(2^16) x^16+x^12+x^3+x+1
GF(2^17) x^17+x^3+1
GF(2^18) x^18+x^7+1
GF(2^19) x^19+x^5+x^2+x+1
GF(2^20) x^20+x^3+1
GF(2^21) x^21+x^2+1
GF(2^22) x^22+x+1
GF(2^23) x^23+x^5+1
GF(2^24) x^24+x^7+x^2+x+1
GF(2^25) x^25+x^3+1
GF(2^26) x^26+x^6+x^2+x+1
GF(2^27) x^27+x^5+x^2+x+1
GF(2^28) x^28+x^3+1
GF(2^29) x^29+x^2+1
GF(2^30) x^30+x^23+x^2+x+1
GF(2^31) x^31+x^3+1
GF(2^32) x^32+x^22+x^2+x+1
GF(2^33) x^33+x^13+1
GF(2^34) x^34+x^8+x^4+x^3+1
GF(2^35) x^35+x^2+1
GF(2^36) x^36+x^11+1
GF(2^37) x^37+x^6+x^4+x+1
GF(2^38) x^38+x^6+x^5+x+1
GF(2^39) x^39+x^4+1
GF(2^40) x^40+x^5+x^4+x^3+1
GF(2^41) x^41+x^3+1
GF(2^42) x^42+x^7+x^4+x^3+1
GF(2^43) x^43+x^6+x^4+x^3+1
GF(2^44) x^44+x^6+x^5+x^2+1
GF(2^45) x^45+x^4+x^3+x+1
GF(2^46) x^46+x^8+x^7+x^6+1
GF(2^47) x^47+x^5+1
GF(2^48) x^48+x^9+x^7+x^4+1
GF(2^49) x^49+x^9+1
GF(2^50) x^50+x^4+x^3+x^2+1
GF(2^51) x^51+x^6+x^3+x+1
GF(2^52) x^52+x^3+1
GF(2^53) x^53+x^6+x^2+x+1
GF(2^54) x^54+x^8+x^6+x^3+1
GF(2^55) x^55+x^24+1
GF(2^56) x^56+x^7+x^4+x^2+1
GF(2^57) x^57+x^7+1
GF(2^58) x^58+x^19+1
GF(2^59) x^59+x^7+x^4+x^2+1
GF(2^60) x^60+x+1
GF(2^61) x^61+x^5+x^2+x+1
GF(2^62) x^62+x^6+x^5+x^3+1
GF(2^63) x^63+x+1
GF(2^64) x^64+x^4+x^3+x+1
GF(2^65) x^65+x^18+1
GF(2^66) x^66+x^9+x^8+x^6+1
GF(2^67) x^67+x^5+x^2+x+1
GF(2^68) x^68+x^9+1
GF(2^69) x^69+x^6+x^5+x^2+1
GF(2^70) x^70+x^5+x^3+x+1
GF(2^71) x^71+x^6+1
GF(2^72) x^72+x^10+x^9+x^3+1
GF(2^73) x^73+x^25+1
GF(2^74) x^74+x^7+x^4+x^3+1
GF(2^75) x^75+x^6+x^3+x+1
GF(2^76) x^76+x^5+x^4+x^2+1
GF(2^77) x^77+x^6+x^5+x^2+1
GF(2^78) x^78+x^7+x^2+x+1
GF(2^79) x^79+x^9+1
GF(2^80) x^80+x^9+x^4+x^2+1
GF(2^81) x^81+x^4+1
GF(2^82) x^82+x^9+x^6+x^4+1
GF(2^83) x^83+x^7+x^4+x^2+1
GF(2^84) x^84+x^13+1
GF(2^85) x^85+x^8+x^2+x+1
GF(2^86) x^86+x^6+x^5+x^2+1
GF(2^87) x^87+x^13+1
GF(2^88) x^88+x^11+x^9+x^8+1
GF(2^89) x^89+x^38+1
GF(2^90) x^90+x^5+x^3+x^2+1
GF(2^91) x^91+x^8+x^5+x+1
GF(2^92) x^92+x^6+x^5+x^2+1
GF(2^93) x^93+x^2+1
GF(2^94) x^94+x^21+1
GF(2^95) x^95+x^11+1
GF(2^96) x^96+x^10+x^9+x^6+1
GF(2^97) x^97+x^6+1
GF(2^98) x^98+x^11+1
GF(2^99) x^99+x^7+x^5+x^4+1
GF(2^100) x^100+x^37+1
GF(2^101) x^101+x^7+x^6+x+1
GF(2^102) x^102+x^6+x^5+x^3+1
GF(2^103) x^103+x^9+1
GF(2^104) x^104+x^11+x^10+x+1
GF(2^105) x^105+x^16+1
GF(2^106) x^106+x^15+1
GF(2^107) x^107+x^9+x^7+x^4+1
GF(2^108) x^108+x^31+1
GF(2^109) x^109+x^5+x^4+x^2+1
GF(2^110) x^110+x^6+x^4+x+1
GF(2^111) x^111+x^10+1
GF(2^112) x^112+x^11+x^6+x^4+1
GF(2^113) x^113+x^9+1
GF(2^114) x^114+x^11+x^2+x+1
GF(2^115) x^115+x^8+x^7+x^5+1
GF(2^116) x^116+x^6+x^5+x^2+1
GF(2^117) x^117+x^5+x^2+x+1
GF(2^118) x^118+x^33+1
GF(2^119) x^119+x^8+1
GF(2^120) x^120+x^9+x^6+x^2+1
GF(2^121) x^121+x^18+1
GF(2^122) x^122+x^6+x^2+x+1
GF(2^123) x^123+x^2+1
GF(2^124) x^124+x^37+1
GF(2^125) x^125+x^7+x^6+x^5+1
GF(2^126) x^126+x^7+x^4+x^2+1
GF(2^127) x^127+x+1
GF(2^128) x^128+x^7+x^2+x+1
GF(2^144) x^144+x^7+x^4+x^2+1
GF(2^160) x^160+x^5+x^3+x^2+1
GF(2^176) x^176+x^12+x^11+x^9+1
GF(2^192) x^192+x^15+x^11+x^5+1
GF(2^200) x^200+x^5+x^3+x^2+1
GF(2^208) x^208+x^9+x^3+x+1
GF(2^224) x^224+x^12+x^7+x^2+1
GF(2^240) x^240+x^8+x^5+x^3+1
GF(2^256) x^256+x^10+x^5+x^2+1
GF(2^300) x^300+x^7+1
GF(2^320) x^320+x^4+x^3+x+1
GF(2^360) x^360+x^26+x^25+x+1
GF(2^384) x^384+x^16+x^15+x^6+1
GF(2^400) x^400+x^5+x^3+x^2+1
GF(2^480) x^480+x^16+x^13+x^7+1
GF(2^512) x^512+x^8+x^5+x^2+1
GF(2^600) x^600+x^11+x^10+x+1
GF(2^720) x^720+x^11+x^8+x^2+1
GF(2^840) x^840+x^11+x^5+x+1
GF(2^960) x^960+x^13+x^9+x^6+1
GF(2^1200) x^1200+x^23+x^8+x^5+1

# Примитивные неприводимые многочлены над полем GF(3)

GF(3^2) x^2+x+2
GF(3^3) x^3+2*x+1
GF(3^4) x^4+x+2
GF(3^5) x^5+2*x+1
GF(3^6) x^6+x+2
GF(3^7) x^7+2*x^2+1
GF(3^8) x^8+x^3+2
GF(3^9) x^9+2*x^4+1
GF(3^10) x^10+x^3+x+2
GF(3^11) x^11+2*x^2+1
GF(3^12) x^12+x^5+x+2
GF(3^13) x^13+2*x+1
GF(3^14) x^14+x+2
GF(3^15) x^15+2*x^2+1
GF(3^16) x^16+x^7+2
GF(3^17) x^17+2*x+1
GF(3^18) x^18+x^9+x^5+2
GF(3^19) x^19+2*x^2+1
GF(3^20) x^20+x^5+x+2
GF(3^21) x^21+2*x^5+1
GF(3^22) x^22+x^5+2
GF(3^23) x^23+2*x^3+1
GF(3^24) x^24+x^13+x^5+2
GF(3^25) x^25+2*x^3+1
GF(3^26) x^26+x^7+2
GF(3^27) x^27+2*x^7+1
GF(3^28) x^28+x^13+2
GF(3^29) x^29+2*x^4+1
GF(3^30) x^30+x+2
GF(3^31) x^31+2*x^5+1
GF(3^32) x^32+x^5+2
GF(3^33) x^33+2*x^5+1
GF(3^34) x^34+x^3+x+2
GF(3^35) x^35+2*x^2+1
GF(3^36) x^36+x^17+x+2
GF(3^37) x^37+2*x^6+1
GF(3^38) x^38+x^13+x^5+2
GF(3^39) x^39+2*x^5+x^4+1
GF(3^40) x^40+x+2
GF(3^41) x^41+2*x+1
GF(3^42) x^42+x^9+x^7+2
GF(3^43) x^43+2*x^17+1
GF(3^44) x^44+x^3+2
GF(3^45) x^45+2*x^17+1
GF(3^46) x^46+x^5+2
GF(3^47) x^47+2*x^15+1
GF(3^48) x^48+x^11+x^6+2*x^4+2
GF(3^49) x^49+x^9+2*x^6+1
GF(3^50) x^50+x^11+x^9+2
GF(3^51) x^51+2*x+1
GF(3^52) x^52+x^7+2
GF(3^53) x^53+2*x^13+1
GF(3^54) x^54+x+2
GF(3^55) x^55+2*x^23+1
GF(3^56) x^56+x^3+2
GF(3^57) x^57+x^7+2*x^2+1
GF(3^58) x^58+x^13+x^11+2
GF(3^59) x^59+2*x^17+1
GF(3^60) x^60+x^5+x+2
GF(3^61) x^61+2*x^7+1
GF(3^62) x^62+x^9+x^7+2
GF(3^63) x^63+2*x^26+1
GF(3^64) x^64+x^3+2
GF(3^72) x^72+x^18+x^3+2*x^2+2
GF(3^80) x^80+x^21+2
GF(3^96) x^96+x^7+x^6+2*x^4+2
GF(3^100) x^100+x^17+x+2
GF(3^112) x^112+x^43+2
GF(3^128) x^128+x^5+2*x^3+x^2+2
GF(3^144) x^144+x^5+2*x^4+x^2+2
GF(3^160) x^160+x^27+2
GF(3^176) x^176+x^15+2
GF(3^192) x^192+x^5+2*x^4+x^2+2
GF(3^200) x^200+x^3+2
GF(3^208) x^208+x^51+2
GF(3^224) x^224+x^23+2
GF(3^240) x^240+x^35+x^19+2
GF(3^256) x^256+x^7+2*x^3+x^2+2
GF(3^300) x^300+x^9+2*x^6+x^4+2

# Примитивные неприводимые многочлены над полем GF(5)

GF(5^2) x^2+x+2
GF(5^3) x^3+3*x+2
GF(5^4) x^4+x^2+2*x+2
GF(5^5) x^5+x^2+2
GF(5^6) x^6+x+2
GF(5^7) x^7+3*x+2
GF(5^8) x^8+x^2+2*x+3
GF(5^9) x^9+2*x^4+3
GF(5^10) x^10+x^2+x+3
GF(5^11) x^11+x^2+2
GF(5^12) x^12+x^3+2*x+3
GF(5^13) x^13+2*x^6+3
GF(5^14) x^14+x^9+x+3
GF(5^15) x^15+x^2+2
GF(5^16) x^16+x^3+3*x+2
GF(5^17) x^17+x^14+2
GF(5^18) x^18+x^4+2*x+2
GF(5^19) x^19+4*x^9+2
GF(5^20) x^20+x^2+2*x+3
GF(5^21) x^21+4*x+2
GF(5^22) x^22+x^5+2
GF(5^23) x^23+2*x^2+3
GF(5^24) x^24+x^3+2*x^2+2
GF(5^25) x^25+3*x^7+2
GF(5^26) x^26+x^5+4*x^3+3
GF(5^27) x^27+4*x+2
GF(5^28) x^28+x^3+2*x+3
GF(5^29) x^29+2*x^6+3
GF(5^30) x^30+x^5+3*x^2+3
GF(5^31) x^31+3*x+2
GF(5^32) x^32+x^5+2*x^3+3
GF(5^36) x^36+x^7+3*x+2
GF(5^40) x^40+x^11+2*x^8+2
GF(5^48) x^48+x^7+4*x^6+3
GF(5^56) x^56+x^7+4*x^6+3
GF(5^64) x^64+x^7+2*x^4+2
GF(5^72) x^72+x^6+2*x^5+2
GF(5^80) x^80+x^5+2*x^2+2
GF(5^96) x^96+x^3+4*x^2+2
GF(5^100) x^100+x^9+3*x^6+3
GF(5^112) x^112+x^7+4*x^2+2
GF(5^128) x^128+x^3+x+3
GF(5^144) x^144+x^15+3*x^10+3
GF(5^160) x^160+x^6+2*x^5+3
GF(5^200) x^200+x^8+x^5+3

# Примитивные неприводимые многочлены над полем GF(7)

GF(7^2) x^2+x+3
GF(7^3) x^3+3*x+2
GF(7^4) x^4+x^2+3*x+5
GF(7^5) x^5+x+4
GF(7^6) x^6+x^3+x+5
GF(7^7) x^7+x^4+2
GF(7^8) x^8+x+3
GF(7^9) x^9+3*x^2+4
GF(7^10) x^10+x^5+x+3
GF(7^11) x^11+x+4
GF(7^12) x^12+x^5+3*x+5
GF(7^13) x^13+5*x^2+2
GF(7^14) x^14+x^9+3
GF(7^15) x^15+x^8+5*x^2+4
GF(7^16) x^16+x^15+3
GF(7^17) x^17+x+4
GF(7^18) x^18+x^7+6*x+3
GF(7^19) x^19+x^8+4
GF(7^20) x^20+x^3+3
GF(7^21) x^21+3*x^8+4
GF(7^22) x^22+x^3+3
GF(7^23) x^23+x^10+4
GF(7^24) x^24+x^5+6*x+3
GF(7^25) x^25+x^4+2
GF(7^26) x^26+x^9+3
GF(7^27) x^27+3*x^8+4
GF(7^28) x^28+x^4+3*x+3
GF(7^29) x^29+x^13+4
GF(7^30) x^30+x^2+x+5
GF(7^31) x^31+x^4+2
GF(7^32) x^32+x^7+3
GF(7^36) x^36+x^5+3*x^3+5
GF(7^40) x^40+x^9+3
GF(7^48) x^48+x^5+3*x+5
GF(7^56) x^56+x^2+x+5
GF(7^64) x^64+x^21+3
GF(7^72) x^72+x^9+x+5
GF(7^80) x^80+x^69+3
GF(7^96) x^96+x^7+x^3+5
GF(7^100) x^100+x^5+5*x+3
GF(7^112) x^112+x^7+5*x^4+3
GF(7^128) x^128+x^6+3*x^3+3
GF(7^144) x^144+x^5+4*x+5
GF(7^160) x^160+x^5+x^4+5
GF(7^200) x^200+x^2+x+3
# Примитивные неприводимые многочлены над полем GF(11)

GF(11^2) x^2+x+7
GF(11^3) x^3+x+4
GF(11^4) x^4+x+2
GF(11^5) x^5+2*x^2+9
GF(11^6) x^6+x^2+2*x+8
GF(11^7) x^7+x+4
GF(11^8) x^8+x^2+2*x+6
GF(11^12) x^12+x+7
GF(11^16) x^16+x^7+7
GF(11^24) x^24+x+2
GF(11^32) x^32+x^11+7
GF(11^48) x^48+x^11+8
GF(11^64) x^64+x^3+8
GF(11^80) x^80+x^4+2*x+8
GF(11^96) x^96+x^8+4*x+8
GF(11^100) x^100+x^3+4*x^2+6

# Примитивные неприводимые многочлены над полем GF(13)

GF(13^2) x^2+x+2
GF(13^3) x^3+x+6
GF(13^4) x^4+x^2+x+2
GF(13^5) x^5+3*x^2+2
GF(13^6) x^6+x^2+2*x+2
GF(13^7) x^7+x^4+2
GF(13^8) x^8+x^3+x+2
GF(13^12) x^12+x^2+x+2
GF(13^16) x^16+x^3+6
GF(13^24) x^24+x^2+6*x+2
GF(13^32) x^32+x^4+2*x+11
GF(13^48) x^48+x^2+2*x+6
GF(13^64) x^64+x^3+x+11
GF(13^80) x^80+x^3+4*x^2+2
GF(13^96) x^96+x^5+8*x^4+6
GF(13^100) x^100+x^4+2*x+2

# Примитивные неприводимые многочлены над полем GF(17)

GF(17^2) x^2+x+3
GF(17^3) x^3+x+3
GF(17^4) x^4+x+11
GF(17^5) x^5+x+3
GF(17^6) x^6+x+12
GF(17^7) x^7+x+5
GF(17^8) x^8+x^3+5
GF(17^12) x^12+x^5+6
GF(17^16) x^16+x^3+2*x+7
GF(17^24) x^24+x^2+2*x+7
GF(17^32) x^32+x^2+x+6
GF(17^48) x^48+x^2+2*x+6
GF(17^64) x^64+x^7+4*x+7
GF(17^80) x^80+x^5+2*x^2+12
GF(17^96) x^96+x^2+8*x+3
GF(17^100) x^100+x^3+x+7

# Примитивные неприводимые многочлены над полем GF(19)

GF(19^2) x^2+x+2
GF(19^3) x^3+x+4
GF(19^4) x^4+2*x+10
GF(19^5) x^5+x+9
GF(19^6) x^6+x+3
GF(19^7) x^7+x^2+6
GF(19^8) x^8+x+2
GF(19^12) x^12+x+15
GF(19^16) x^16+x^2+5*x+13
GF(19^24) x^24+x^5+14
GF(19^32) x^32+x^13+3
GF(19^48) x^48+x^5+2*x+13
GF(19^64) x^64+x^13+2
GF(19^80) x^80+x+14
GF(19^96) x^96+x^4+5*x+13
GF(19^100) x^100+x^2+8*x+3

# Примитивные неприводимые многочлены над полем GF(23)

GF(23^2) x^2+x+7
GF(23^3) x^3+x+3
GF(23^4) x^4+x+11
GF(23^5) x^5+x+3
GF(23^6) x^6+x^5+7
GF(23^7) x^7+x^2+3
GF(23^8) x^8+x^3+7
GF(23^12) x^12+x^5+11
GF(23^16) x^16+x^15+11
GF(23^24) x^24+x+7
GF(23^32) x^32+x^9+19
GF(23^48) x^48+2*x^13+19
GF(23^64) x^64+x^13+11
GF(23^80) x^80+x^33+17

# Примитивные неприводимые многочлены над полем GF(29)

GF(29^2) x^2+x+3
GF(29^3) x^3+x+11
GF(29^4) x^4+x+19
GF(29^5) x^5+x+8
GF(29^6) x^6+x+3
GF(29^7) x^7+x+11
GF(29^8) x^8+x^2+3*x+3
GF(29^12) x^12+x+15
GF(29^16) x^16+x^3+21
GF(29^24) x^24+x+21
GF(29^32) x^32+x+19
GF(29^48) x^48+x^19+19
GF(29^64) x^64+2*x^17+8
GF(29^80) x^80+x^2+x+2

# Примитивные неприводимые многочлены над полем GF(31)

GF(31^2) x^2+x+2
GF(31^3) x^3+x+14
GF(31^4) x^4+x^3+13
GF(31^5) x^5+x+18
GF(31^6) x^6+x^5+12
GF(31^7) x^7+x^2+7
GF(31^8) x^8+x+22
GF(31^12) x^12+x^3+2*x+13
GF(31^16) x^16+x^3+12
GF(31^24) x^24+x^11+22
GF(31^32) x^32+x+12
GF(31^48) x^48+x^35+11
GF(31^64) x^64+x^5+3
GF(31^80) x^80+x^3+12

# Примитивные неприводимые многочлены над полем GF(37)

GF(37^2) x^2+x+5
GF(37^3) x^3+x+13
GF(37^4) x^4+x+2
GF(37^5) x^5+x+5
GF(37^6) x^6+x+20
GF(37^7) x^7+x^2+19
GF(37^8) x^8+x+18
GF(37^12) x^12+x+15
GF(37^16) x^16+x^3+15
GF(37^24) x^24+x^11+18
GF(37^32) x^32+x^17+18
GF(37^48) x^48+x^11+20
GF(37^64) x^64+x^29+22

# Примитивные неприводимые многочлены над полем GF(41)

GF(41^2) x^2+x+12
GF(41^3) x^3+x+6
GF(41^4) x^4+x+17
GF(41^5) x^5+x^3+7
GF(41^6) x^6+x+7
GF(41^7) x^7+x^2+7
GF(41^8) x^8+x^3+15
GF(41^12) x^12+x^3+2*x+12
GF(41^16) x^16+x^7+7
GF(41^24) x^24+x+29
GF(41^32) x^32+x^5+2*x+17
GF(41^48) x^48+x^11+22

# Примитивные неприводимые многочлены над полем GF(43)

GF(43^2) x^2+x+3
GF(43^3) x^3+x+14
GF(43^4) x^4+x+20
GF(43^5) x^5+x+13
GF(43^6) x^6+x^5+3
GF(43^7) x^7+x+9
GF(43^8) x^8+x^3+28
GF(43^12) x^12+x+33
GF(43^16) x^16+x^5+34
GF(43^24) x^24+x^3+x+19
GF(43^32) x^32+x^17+5
GF(43^48) x^48+x+29

# Примитивные неприводимые многочлены над полем GF(47)

GF(47^2) x^2+x+13
GF(47^3) x^3+x+4
GF(47^4) x^4+x+39
GF(47^5) x^5+x+3
GF(47^6) x^6+x+5
GF(47^7) x^7+x+3
GF(47^8) x^8+x+20
GF(47^12) x^12+x^7+22
GF(47^16) x^16+x^5+11
GF(47^24) x^24+x^19+20
GF(47^32) x^32+x^15+30
GF(47^48) x^48+x+20
GF(47^64) x^64+x^13+29

# Примитивные неприводимые многочлены над полем GF(53)

GF(53^2) x^2+x+5
GF(53^3) x^3+x+5
GF(53^4) x^4+x+18
GF(53^5) x^5+x+26
GF(53^6) x^6+x+8
GF(53^7) x^7+x+5
GF(53^8) x^8+x^5+21
GF(53^12) x^12+x+12
GF(53^16) x^16+x+8
GF(53^24) x^24+x^11+2
GF(53^32) x^32+x+27
GF(53^48) x^48+x^2+x+3

# Примитивные неприводимые многочлены над полем GF(59)

GF(59^2) x^2+x+2
GF(59^3) x^3+x+3
GF(59^4) x^4+x+14
GF(59^5) x^5+x+12
GF(59^6) x^6+x+23
GF(59^7) x^7+x+9
GF(59^8) x^8+x+14
GF(59^12) x^12+x+10
GF(59^16) x^16+x+31
GF(59^24) x^24+x+8
GF(59^32) x^32+x^5+55
GF(59^48) x^48+x^11+43

# Примитивные неприводимые многочлены над полем GF(61)

GF(61^2) x^2+x+2
GF(61^3) x^3+x+17
GF(61^4) x^4+x+2
GF(61^5) x^5+x+7
GF(61^6) x^6+x^5+6
GF(61^7) x^7+x^2+10
GF(61^8) x^8+x^3+2
GF(61^12) x^12+x^11+6
GF(61^16) x^16+x+2
GF(61^24) x^24+x^19+2
GF(61^32) x^32+x+17
GF(61^48) x^48+x^17+35
GF(61^64) x^64+4*x+7

# Примитивные неприводимые многочлены над полем GF(67)

GF(67^2) x^2+x+12
GF(67^3) x^3+x+6
GF(67^4) x^4+x+2
GF(67^5) x^5+x+16
GF(67^6) x^6+x^3+x+32
GF(67^7) x^7+x+17
GF(67^8) x^8+x^3+18
GF(67^12) x^12+x^11+18
GF(67^16) x^16+x+28
GF(67^24) x^24+x^7+12
GF(67^32) x^32+x^15+11
GF(67^48) x^48+x^17+32
GF(67^64) x^64+x^3+46

# Примитивные неприводимые многочлены над полем GF(71)

GF(71^2) x^2+x+11
GF(71^3) x^3+x+8
GF(71^4) x^4+x+11
GF(71^5) x^5+x^2+4
GF(71^6) x^6+2*x+13
GF(71^7) x^7+x+4
GF(71^8) x^8+x^3+22
GF(71^12) x^12+2*x+13
GF(71^16) x^16+x^3+47
GF(71^24) x^24+x+56
GF(71^32) x^32+x+11
GF(71^48) x^48+x^5+56

# Примитивные неприводимые многочлены над полем GF(73)

GF(73^2) x^2+x+11
GF(73^3) x^3+x+13
GF(73^4) x^4+x+13
GF(73^5) x^5+x^2+13
GF(73^6) x^6+x+5
GF(73^7) x^7+x^2+13
GF(73^8) x^8+x^3+53
GF(73^12) x^12+x+29
GF(73^16) x^16+x^13+14
GF(73^24) x^24+x^5+15
GF(73^32) x^32+x+47
GF(73^48) x^48+x^3+x+34

# Примитивные неприводимые многочлены над полем GF(79)

GF(79^2) x^2+x+3
GF(79^3) x^3+x+9
GF(79^4) x^4+x+3
GF(79^5) x^5+x^2+4
GF(79^6) x^6+x+6
GF(79^7) x^7+x+4
GF(79^8) x^8+x^3+6
GF(79^12) x^12+x+48
GF(79^16) x^16+x^5+3
GF(79^24) x^24+x^13+30
GF(79^32) x^32+x^9+37
GF(79^48) x^48+x^7+68

# Примитивные неприводимые многочлены над полем GF(83)

GF(83^2) x^2+x+2
GF(83^3) x^3+x+7
GF(83^4) x^4+x+22
GF(83^5) x^5+x+12
GF(83^6) x^6+x+34
GF(83^7) x^7+x^3+10
GF(83^8) x^8+x+8
GF(83^12) x^12+x^5+13
GF(83^16) x^16+x^3+24
GF(83^24) x^24+x^2+x+22
GF(83^32) x^32+x^13+19
GF(83^48) x^48+x+53

# Примитивные неприводимые многочлены над полем GF(89)

GF(89^2) x^2+x+6
GF(89^3) x^3+x+19
GF(89^4) x^4+x+27
GF(89^5) x^5+x+3
GF(89^6) x^6+x+6
GF(89^7) x^7+x^2+15
GF(89^8) x^8+x^5+24
GF(89^12) x^12+x^7+6
GF(89^16) x^16+x^3+15
GF(89^24) x^24+x^11+15
GF(89^32) x^32+x^3+3
GF(89^48) x^48+x^7+28

# Примитивные неприводимые многочлены над полем GF(97)

GF(97^2) x^2+x+5
GF(97^3) x^3+x+7
GF(97^4) x^4+x+23
GF(97^5) x^5+x+7
GF(97^6) x^6+x+10
GF(97^7) x^7+x+13
GF(97^8) x^8+x^5+5
GF(97^12) x^12+x+68
GF(97^16) x^16+x^5+10
GF(97^24) x^24+x+83
GF(97^32) x^32+x^3+5
GF(97^48) x^48+x^11+13 