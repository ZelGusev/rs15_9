/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : Алгоритм Евклида НОД 
--                     поиск НОД
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/
module evklid_nod(
    clk,            // синхросигнал
    rst_n,          // сброс
    en,             // готовность входных данных
    data_i,         // число
    gf,             // поле
    rdy,            // готовность
    data_o          // обратное число
    );
    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    parameter DATA_WIDTH            = 6;
    parameter RAM_WIDTH             = 6;
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input                               clk;            // синхросигнал
    input                               rst_n;          // сброс
    input                               en;             // готовность входных данных
    input    [DATA_WIDTH - 1 : 0]       data_i;         // шина синдрома
    input    [DATA_WIDTH - 1 : 0]       gf;             // поле
    output  reg                         rdy;            // готовность
    output   [DATA_WIDTH - 1 : 0]       data_o;         // шина полином ошибки
    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    reg en_reg;
    reg start;
    integer i;
    integer reg_y;
    integer reg_x;
    reg [DATA_WIDTH - 1 : 0]    reg_gf;
    reg [DATA_WIDTH - 1 : 0]    reg_a;
    reg [DATA_WIDTH - 1 : 0]    reg_b;
    reg [DATA_WIDTH - 1 : 0]    reg_o;
    reg [DATA_WIDTH - 1 : 0]    reg_ab     [RAM_WIDTH];
    //----------------------------------------------------------------------//
    // wires                                                                //
    //----------------------------------------------------------------------//

    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    assign data_o = reg_y;
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//
    always @(posedge clk)
        begin
            if (~rst_n)
                begin
                    en_reg  <= 1'b0;
                    start   <= 1'b0;
                    i <= 0;
                    reg_x   <= 0;
                    reg_y   <= 1;
                    reg_gf  <= 0;
                end
            else
                begin
                    en_reg <= en;
                    if (~en_reg && en)
                        begin
                            reg_y       <= 1;
                            reg_gf      <= gf;
                            reg_ab  [0] <= gf/data_i;
                            reg_a       <= data_i;
                            reg_b       <= gf%data_i;
                            start       <= 1'b1;
                            rdy         <= 1'b0;
                            i           <= i + 1;
                        end
                    else if (start)
                        begin
                            if (reg_a%reg_b != 0)
                                begin
                                    i           <= i + 1;
                                    reg_ab[i]   <= reg_a/reg_b;
                                    reg_a       <= reg_b;
                                    reg_b       <= reg_a%reg_b;
                                end
                            else
                                begin
                                    if (i != 0)
                                        begin
                                            reg_y   <= reg_x - reg_y*reg_ab[i - 1];
                                            reg_x   <= reg_y;
                                            i       <= i - 1;
                                        end
                                    else
                                        begin
                                            rdy     <= 1'b1;
                                            start   <= 1'b0;
                                            i <= 0;
                                            reg_x   <= 0;
                                            reg_gf  <= 0;
                                            if (reg_y < 0)
                                                begin
                                                    reg_y   <= reg_gf + reg_y;
                                                end
                                        end
                                end
                        end
                end
        end
endmodule