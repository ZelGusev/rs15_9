/*************************************************************************************************************
--    Система        : 
--    Разработчик    :
--    Автор          : Гусев Игорь
--
--    Назначение     : Этот пакет (package) содержит компоненты среды тестового окружения
-—                     
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/
`ifndef _GUARD_ENV_PKG_
    `define _GUARD_ENV_PKG_

package tb_env_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tb_scoreboard.svh"
    `include "tb_env.svh"
      
endpackage : tb_env_pkg

`endif // _GUARD_ENV_PKG_