/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : Умножение в поле Галуа 2**3
--                     Производит умножение, затем деление на порождающий полином x**4 + x + 1
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/
module gf2_3mult(
    data_a,         // шина данных
    data_b,         // шина данных
    data_out        // шина результирующих данных
    );
    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    localparam DATA_WIDTH           = 4;
    localparam DATA_MULT_WIDTH      = 7;
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input    [DATA_WIDTH - 1 : 0]       data_a;         // шина данных
    input    [DATA_WIDTH - 1 : 0]       data_b;         // шина данных
    output   [DATA_WIDTH - 1 : 0]       data_out;       // шина результирующих данных
    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // wires                                                                //
    //----------------------------------------------------------------------//
    wire    [DATA_MULT_WIDTH - 1 : 0]   mult;
    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    // умножение
    assign mult[0]  = (data_a[0] & data_b[0]);
    assign mult[1]  = (data_a[0] & data_b[1]) ^ (data_a[1] & data_b[0]);
    assign mult[2]  = (data_a[0] & data_b[2]) ^ (data_a[1] & data_b[1]) ^ (data_a[2] & data_b[0]);
    assign mult[3]  = (data_a[0] & data_b[3]) ^ (data_a[1] & data_b[2]) ^ (data_a[2] & data_b[1]) ^ (data_a[3] & data_b[0]);
    assign mult[4]  = (data_a[1] & data_b[3]) ^ (data_a[2] & data_b[2]) ^ (data_a[3] & data_b[1]);
    assign mult[5]  = (data_a[2] & data_b[3]) ^ (data_a[3] & data_b[2]);
    assign mult[6]  = (data_a[3] & data_b[3]);

    // остаток от деления на порождающий полином x**4 + x + 1
    assign data_out[0] = mult[0] ^ mult[4];
    assign data_out[1] = mult[1] ^ mult[4] ^ mult[5];
    assign data_out[2] = mult[2] ^ mult[5] ^ mult[6];
    assign data_out[3] = mult[3] ^ mult[6];
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//

endmodule