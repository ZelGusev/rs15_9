/*************************************************************************************************************
--    Система        : 
--    Разработчик    : 
--    Автор          : Гусев Игорь
--
--    Назначение     : Сумматор в поле Галуа
--                     Считает сумму в поле обычный xor
--------------------------------------------------------------------------------------------------------------
--    Примечание     : 
*************************************************************************************************************/
module gf2_add(
    data_a,         // шина данных
    data_b,         // шина данных
    data_out        // шина результирующих данных
    );
    //----------------------------------------------------------------------//
    // external parameters                                                  //
    //----------------------------------------------------------------------//
    parameter DATA_WIDTH            = 4;
    //----------------------------------------------------------------------//
    // internal parameters                                                  //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // external signals                                                     //
    //----------------------------------------------------------------------//
    input    [DATA_WIDTH - 1 : 0]       data_a;         // шина данных
    input    [DATA_WIDTH - 1 : 0]       data_b;         // шина данных
    output   [DATA_WIDTH - 1 : 0]       data_out;       // шина результирующих данных
    //----------------------------------------------------------------------//
    // registers                                                            //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // wires                                                                //
    //----------------------------------------------------------------------//
    //----------------------------------------------------------------------//
    // assigns                                                              //
    //----------------------------------------------------------------------//
    // сумматор в поле Галуа
    assign data_out = data_a ^ data_b;
    //----------------------------------------------------------------------//
    // logic                                                                //
    //----------------------------------------------------------------------//

endmodule